/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/mem_group_share/mem.sv