module wta_1
#(parameter NUM_INPUTS = 16)
(
    input logic rst,
    input logic [NUM_INPUTS-1:0] input_spikes,
    output logic [NUM_INPUTS-1:0] output_spikes
);



endmodule: wta_1