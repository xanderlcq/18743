/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/mux_b_t_s/mux_b_t_s.sv