/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/mux/mux.sv