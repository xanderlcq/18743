/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/mux_t_be_t_N/mux_t_be_t_N.sv