/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/lib/sr_latch.sv