/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/mux_b_t_t_n/mux_b_t_t_n.sv