/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/binary2unary/binary2unary.sv