/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/snl/neuron_snl_grl.sv