/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/less_than_eq/less_than_eq.sv