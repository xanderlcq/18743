/afs/andrew.cmu.edu/usr24/sganiger/private/18743/project/18743/src/rtl/greater_than_eq/greater_than_eq.sv