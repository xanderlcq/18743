/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/mem/mem.sv