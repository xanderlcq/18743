/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/wta_1/wta_1.sv