/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/kwta/kwta.sv