/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/wta_1/wrapper.sv