/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/greater_than_eq/greater_than_eq.sv