/afs/andrew.cmu.edu/usr4/kbhat2/private/18-743/project/src/rtl/exclusive_max/exclusive_max.sv