/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/naive_delay/naive_delay.sv