/afs/andrew.cmu.edu/usr24/sganiger/private/18743/project/18743/src/rtl/less_than_eq/less_than_eq.sv