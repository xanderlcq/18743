module tb();

endmodule