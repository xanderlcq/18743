/afs/ece.cmu.edu/usr/acli/Private/18743/src/rtl/kwta_no_tie_break/kwta_no_tie_break.sv